module NOT_gate(
    input   A,
    output  Y_not
);

    assign Y_not = ~A;

endmodule