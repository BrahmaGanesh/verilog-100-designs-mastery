module XOR_gate(
    input   A,
    input   B,
    output  Y_xor
);

    assign Y_xor = A ^ B;

endmodule