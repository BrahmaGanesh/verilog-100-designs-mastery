module AND_gate(
    input   A,
    input   B,
    output  Y_and
);

    assign Y_and = A & B;

endmodule