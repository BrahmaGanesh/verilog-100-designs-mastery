module buffer(
    input   A,
    output  Y_buff
);

    assign Y_buff = A;

endmodule